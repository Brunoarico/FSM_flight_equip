LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY selector IS
	PORT (
		SEL : STD_LOGIC_VECTOR(1 DOWNTO 0);
		D0A : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		D1A : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		D2A : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		D3A : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		D0T : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		D1T : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		D2T : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		D3T : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		D0P : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		D1P : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		D2P : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		D3P : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		D0C : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		D1C : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		D2C : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		D3C : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		D0 : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		D1 : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		D2 : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		D3 : OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
	);
END selector;

ARCHITECTURE Behavioral OF selector IS

BEGIN
	PROCESS (SEL)
	BEGIN
		IF SEL = "00" THEN
			D0 <= D0C;
			D1 <= D1C;
			D2 <= D2C;
			D3 <= D3C;
		ELSIF SEL = "01" THEN
			D0 <= D0T;
			D1 <= D1T;
			D2 <= D2T;
			D3 <= D3T;
		ELSIF SEL = "10" THEN
			D0 <= D0A;
			D1 <= D1A;
			D2 <= D2A;
			D3 <= D3A;
		ELSIF SEL = "11" THEN
			D0 <= D0P;
			D1 <= D1P;
			D2 <= D2P;
			D3 <= D3P;
		END IF;
	END PROCESS;

END Behavioral;