LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY bcd_converter IS
	PORT (
		BIN : IN STD_LOGIC_VECTOR(3 DOWNTO 0); -- Entrada BCD de 4 bits
		SEGS : OUT STD_LOGIC_VECTOR(6 DOWNTO 0) -- Saída para os segmentos do display de 7 segmentos
	);
END bcd_converter;

ARCHITECTURE Behavioral OF bcd_converter IS
BEGIN
	SEGS <= "1000000" WHEN BIN = "0000" ELSE -- 0
		"1111001" WHEN BIN = "0001" ELSE -- 1
		"0100100" WHEN BIN = "0010" ELSE -- 2 
		"0110000" WHEN BIN = "0011" ELSE -- 3
		"0011001" WHEN BIN = "0100" ELSE -- 4
		"0010010" WHEN BIN = "0101" ELSE -- 5
		"0000010" WHEN BIN = "0110" ELSE -- 6
		"1111000" WHEN BIN = "0111" ELSE -- 7
		"0000000" WHEN BIN = "1000" ELSE -- 8
		"0011000" WHEN BIN = "1001" ELSE -- 9
		"0111111" WHEN BIN = "1010" ELSE -- -
		"0111000" WHEN BIN = "1011" ELSE -- L
		"1000110" WHEN BIN = "1100" ELSE -- C
		"1111111" WHEN BIN = "1101" ELSE -- Desligado
		"0001000" WHEN BIN = "1110" ELSE -- A
		"0001100" WHEN BIN = "1111" ELSE -- F
		"0000000";
END Behavioral;